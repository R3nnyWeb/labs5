module v82 (c,q,y);
input c;
output [2:0]q;
output [2:0] y;
reg [2:0] q;
always @ (posedge c) if (q  == 7) q = 2; else q = q + 1;
assign y[2] = ~q[2] & q[1] & ~q[0] | q[2] & q[1] & ~q[0] | q[2]& q[1] & q[0];
assign y[1] = q[2] & ~q[1] & ~q[0] | q[2] & ~q[1] & q[0] | q[2]& q[1] & ~q[0];
assign y[0] = ~q[2] & q[1] & ~q[0] | ~q[2] & q[1] & q[0] | q[2]& ~q[1] & ~q[0];
endmodule